`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: University of Thessaly
// Engineer: Dimitris Voitsidis
// 
// Create Date: 12/08/2023 11:07:23 AM
// Design Name: Counter
// Module Name: counter
// Project Name: Universal Asynchronous Receiver Transmitter — UART
// Target Devices: Artix 7
// Tool Versions: 
// Description: A parameterized, for size, counter with hold.
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
///////////////////////////////////////////////////////////////////////////////////////////////////


module counter #(parameter size=8) (reset, clk, hold, counter);
  input reset, clk, hold;
  output reg [size-1:0] counter;

  always @ (posedge clk or posedge reset)
  begin
    if(reset)
    begin
      counter <= 0;
    end
    else
    if(hold)
    begin
      counter <= counter;
    end
    else
    begin
      counter <= counter + 1'b1;
    end 
  end
endmodule